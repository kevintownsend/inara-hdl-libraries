module switch_8_8(clk, rst, p0_push_in, p0_route, p0_stall_in, p0_push_out, p0_stall_out,/* TODO the rest */);

endmodule
