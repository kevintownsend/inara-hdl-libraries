module linked_fifo(rst, clk, push, push_fifo, pop, pop_fifo, d, q, empty, full, count);
    parameter WIDTH = 8;
    parameter DEPTH = 32;
    parameter FIFOS = 8;
    parameter FIFO_LOG2 = 3
    parameter DEPTH_LOG2 = 0;
    //TODO finish
endmodule
