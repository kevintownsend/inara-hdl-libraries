function integer abs;
    input integer value;
    if (value < 0)
        abs=-value;
    else
        abs=value;
endfunction
