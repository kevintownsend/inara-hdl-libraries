`define DEBUG 0
